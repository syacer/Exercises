library verilog;
use verilog.vl_types.all;
entity TestAddSub1Bit is
end TestAddSub1Bit;
